/*-
 * Copyright (c) 2018 Krzysztof Piotr Koch
 * All rights reserved.
 *
 * Redistribution and use in source and binary forms, with or without
 * modification, are permitted provided that the following conditions
 * are met:
 * 1. Redistributions of source code must retain the above copyright
 *    notice, this list of conditions and the following disclaimer.
 * 2. Redistributions in binary form must reproduce the above copyright
 *    notice, this list of conditions and the following disclaimer in the
 *    documentation and/or other materials provided with the distribution.
 *
 * THIS SOFTWARE IS PROVIDED BY THE AUTHOR AND CONTRIBUTORS ``AS IS'' AND
 * ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
 * IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
 * ARE DISCLAIMED.  IN NO EVENT SHALL THE AUTHOR OR CONTRIBUTORS BE LIABLE
 * FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
 * DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
 * OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
 * HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
 * LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
 * OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
 * SUCH DAMAGE.
 */


/*-
 * Instrution decoder for every instruction in RV32IM and RV64IM 
 * (user-level ISA)
 */

// ------------------------------------------------------------------------
// Instruction decoder
// ------------------------------------------------------------------------
function Action instr_decode(Instr instr);
    action
        case (instr) matches
// ----------------------------------------------------------------------------
// RV32I Base Instruction Set 
// ----------------------------------------------------------------------------
            
            // I-type (jalr) 
            //  ____________________________________
            // |  imm[11:0] | rs1 | f3|  rd | opcode|
            32'b????????????_?????_000_?????_1100111:   jalr(instr);
            32'b????????????_?????_000_?????_0010011:   addi(instr);
            32'b????????????_?????_010_?????_0010011:   slti(instr);
            32'b????????????_?????_011_?????_0010011:   sltiu(instr);
            32'b????????????_?????_100_?????_0010011:   xori(instr);
            32'b????????????_?????_110_?????_0010011:   ori(instr);
            32'b????????????_?????_111_?????_0010011:   andi(instr);
            32'b????????????_?????_000_?????_0000011:   lb(instr);
            32'b????????????_?????_001_?????_0000011:   lh(instr);
            32'b????????????_?????_010_?????_0000011:   lw(instr);
            32'b????????????_?????_100_?????_0000011:   lbu(instr);
            32'b????????????_?????_101_?????_0000011:   lhu(instr);

            // I-type (shifts)
`ifdef RV32 
            // RV32
            //  _____________________________________
            // | func7 |shamt| rs1 | f3|  rd | opcode|
            32'b0000000_?????_?????_001_?????_0010011:  slli(instr);
            32'b0000000_?????_?????_101_?????_0010011:  srli(instr);
            32'b0100000_?????_?????_101_?????_0010011:  srai(instr);
`elsif RV64
            // RV64
            //  _____________________________________
            // |      | shamt| rs1 | f3|  rd | opcode|
            32'b000000_??????_?????_001_?????_0010011:  slli(instr);
            32'b000000_??????_?????_101_?????_0010011:  srli(instr);
            32'b010000_??????_?????_101_?????_0010011:  srai(instr);
`endif
            // B-type
            //  _________________________________________________
            // |imm[12|10:5]| rs2 | rs1 | f3| imm[4:1|11]| opcode|
            32'b____?_??????_?????_?????_000_______????_?_1100011:  beq(instr);
            32'b____?_??????_?????_?????_001_______????_?_1100011:  bne(instr);
            32'b____?_??????_?????_?????_100_______????_?_1100011:  blt(instr);
            32'b____?_??????_?????_?????_101_______????_?_1100011:  bge(instr);
            32'b____?_??????_?????_?????_110_______????_?_1100011:  bltu(instr);
            32'b____?_??????_?????_?????_111_______????_?_1100011:  bgeu(instr);
            
            // S-type
            //  ___________________________________________
            // | imm[11:5]| rs2 | rs1 | f3|imm[4:0]| opcode|
            32'b___???????_?????_?????_000____?????_0100011:    sb(instr);
            32'b___???????_?????_?????_001____?????_0100011:    sh(instr);
            32'b___???????_?????_?????_010____?????_0100011:    sw(instr);
 
            // R-type
            //  _____________________________________
            // | func7 | rs2 | rs1 | f3|  rd | opcode|
            32'b0000000_?????_?????_000_?????_0110011:  addR(instr);
            32'b0100000_?????_?????_000_?????_0110011:  subR(instr);
            32'b0000000_?????_?????_001_?????_0110011:  sllR(instr);
            32'b0000000_?????_?????_010_?????_0110011:  sltR(instr);
            32'b0000000_?????_?????_011_?????_0110011:  sltuR(instr);
            32'b0000000_?????_?????_100_?????_0110011:  xorR(instr);
            32'b0000000_?????_?????_101_?????_0110011:  srlR(instr);
            32'b0100000_?????_?????_101_?????_0110011:  sraR(instr);
            32'b0000000_?????_?????_110_?????_0110011:  orR(instr);
            32'b0000000_?????_?????_111_?????_0110011:  andR(instr);

            // MISC-MEM instructions
            //  ______________________________________
            // |    |pred|succ| rs1 | f3|  rd | opcode|
            32'b0000_????_????_00000_000_00000_0001111: fence(instr);
            32'b0000_0000_0000_00000_001_00000_0001111: fencei(instr);

            // Environment Call and Breakpoints
            //  ____________________________________
            // |            | rs1 | f3|  rd | opcode|
            32'b000000000000_00000_000_00000_1110011:   ecall(instr);
            32'b000000000001_00000_000_00000_1110011:   ebreak(instr);

            // Systen Instructions
            //  ____________________________________
            // |     csr    | rs1 | f3|  rd | opcode|
            32'b????????????_?????_001_?????_1110011:   csrrw(instr);
            32'b????????????_?????_010_?????_1110011:   csrrs(instr);
            32'b????????????_?????_011_?????_1110011:   csrrc(instr);
            //  ____________________________________
            // |     csr    | zimm| f3|  rd | opcode|
            32'b????????????_?????_101_?????_1110011:   csrrwi(instr);
            32'b????????????_?????_110_?????_1110011:   csrrsi(instr);
            32'b????????????_?????_111_?????_1110011:   csrrci(instr);
`ifdef RVxxM
// ----------------------------------------------------------------------------
// RV32M Standard Extension (multiply and divide)
// ----------------------------------------------------------------------------
            // R-type
            //  _____________________________________
            // | func7 | rs2 | rs1 | f3|  rd | opcode|       
            32'b0000001_?????_?????_000_?????_0110011:  mul(instr); 
            32'b0000001_?????_?????_001_?????_0110011:  mulh(instr);            
            32'b0000001_?????_?????_010_?????_0110011:  mulhsu(instr);            
            32'b0000001_?????_?????_011_?????_0110011:  mulhu(instr);            
            32'b0000001_?????_?????_100_?????_0110011:  div(instr);            
            32'b0000001_?????_?????_101_?????_0110011:  divu(instr);            
            32'b0000001_?????_?????_110_?????_0110011:  rem(instr);            
            32'b0000001_?????_?????_111_?????_0110011:  remu(instr);            
`endif              

`ifdef RV64 
// ----------------------------------------------------------------------------
// RV64I Base Instruction Set (in addition to RV32I)
// ----------------------------------------------------------------------------
            // I-type
            //  ____________________________________
            // |  imm[11:0] | rs1 | f3|  rd | opcode|
            32'b????????????_?????_000_?????_0011011:   addiw(instr);

            // I-type (shifts)
            //  _____________________________________
            // | func7 |shamt| rs1 | f3|  rd | opcode|
            32'b0000000_?????_?????_001_?????_0011011:  slliw(instr);
            32'b0000000_?????_?????_101_?????_0011011:  srliw(instr);
            32'b0100000_?????_?????_101_?????_0011011:  sraiw(instr);

            // R-type
            //  _____________________________________
            // | func7 | rs2 | rs1 | f3|  rd | opcode|
            32'b0000000_?????_?????_000_?????_0111011:  addw(instr);
            32'b0100000_?????_?????_000_?????_0111011:  subw(instr);
            32'b0000000_?????_?????_001_?????_0111011:  sllw(instr);
            32'b0000000_?????_?????_101_?????_0111011:  srlw(instr);
            32'b0100000_?????_?????_101_?????_0111011:  sraw(instr);
`endif
            
            // J-type
            //  _____________________________________
            // | imm[20|10:1|11|19:12] |  rd | opcode|
            32'b?_?????????_?_?????????_?????_1101111:  jal(instr);

            // U-type
            //  __________________________________
            // |     imm[31:13]     |  rd | opcode|
            32'b????????????????????_?????_0110111:     lui(instr);
            32'b????????????????????_?????_0010111:     auipc(instr);

            default: raiseException(EXC_ILLEGAL_INSTR, pc.read(), 
                                    tagged Fault_Instr instr);
        endcase
    endaction
endfunction

